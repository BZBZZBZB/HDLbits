module top_module (
    input clk,
    input areset,
    input x,
    output z
); 

endmodule